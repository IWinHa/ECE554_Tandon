module MAC #(parameter DATA_WIDTH = 8) (
	input clk,
	input rst_n,
	input En,
	input Clr,
	input [DATA_WIDTH-1:0] Ain,
	input [DATA_WIDTH-1:0] Bin,
	output reg [DATA_WIDTH*3-1:0] Cout
);


always_ff @(posedge clk or negedge rst_n) begin
	if (~rst_n) Cout <= {(DATA_WIDTH*3-1){1'b0}};
	else if (Clr) Cout <= {(DATA_WIDTH*3-1){1'b0}};
	else if (En) Cout <= (Ain * Bin) + Cout;
end
	

endmodule
